package clk_pkg;
    `include "cfg_clk.sv"
    `include "driver_clk.sv"
    `include "agent_clk.sv"
endpackage : clk_pkg
