package rst_pkg;
    `include "transaction_reset.sv"
    `include "driver_reset.sv"
    `include "sequencer_reset.sv"
    `include "seq_reset.sv"
    `include "agent_reset.sv"
endpackage : rst_pkg
