`include "base_test.sv"

//testcases:
`include "test_i2c_write.sv"
`include "test_i2c_read.sv"

`include "test_adc_read.sv"

`include "test_regs_ral.sv"

`include "test_dummy.sv"

`include "test_fir.sv"
`include "test_cic.sv"

`include "test_reset.sv"
