package i2c_pkg;
    `include "cfg_i2c.sv"
    `include "transaction_i2c.sv"
    `include "monitor_i2c.sv"
    `include "driver_i2c.sv"
    `include "seq_i2c.sv"
    `include "agent_i2c.sv"
    `include "adapter_i2c.sv"
endpackage : i2c_pkg
